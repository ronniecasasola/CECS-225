`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:16:00 10/24/2016 
// Design Name: 
// Module Name:    flopr 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module flopr(
    input clk,
    input reset,
    input [7:0] d,
    output reg [7:0] q
    );

always @(posedge clk, posedge reset)
	if( reset ) q = 0;
	else			q = d;

endmodule
