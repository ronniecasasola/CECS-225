`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:26:05 10/24/2016 
// Design Name: 
// Module Name:    datapath 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module datapath(
    input clk,
    input reset,
    input memtoreg,
    input pcsrc,
    input alusrc,
    input regdst,
    input regwrite,
    input jump,
    input [2:0] alucontrol,
    input [31:0] instr,
    input [31:0] readdata,
    output zero,
    output [31:0] pc,
    output [31:0] aluresult,
    output [31:0] writedata
    );

wire [4:0] writereg;
wire [31:0] pcnext, pcnextbr, pcplus4, pcbranch;
wire [31:0] signimm, signimmsh;
wire [31:0] srca, srcb, result;
/**************** next PC logic **************/
//program counter
flopr		pcreg(	.clk(	clk			),
						.reset(	reset		),
						.d(	pcnext[7:0]),
						.q(	pc[7:0]		));
						
//Adder to increment the PC value
Adder_32 pcadd1(	.augend(	pc	),
						.addend( 32'h4 ),
						.sum(	pcplus4 ));
						
// shift left the sign extended constant
sl2	immsh(	.a(	signimm		),
					.y(	signimmsh	));
						
//branch address adder
Adder_32 pcadd2(	.augend(	signimmsh	),
						.addend(	pcplus4		),
						.sum(	pcbranch		));
						
//branch mux
mux2_32 pcbrmux(	.in0(	pcplus4	),
						.in1(	pcbranch	),
						.sel(	pcsrc		),
						.out(	pcnextbr	));
						
//jump mux
mux2_32 pcmux(		.in0(	pcnextbr	),
						.in1( {pcplus4[31:28], instr[25:0], 2'b00}),
						.sel(	jump		),
						.out(	pcnext	));

/****************************************/

/****************** register file logic************/
// The register file
regfile rf(			.clk(	clk		),
						.we3(	regwrite	),
						.ra1(	instr[25:21]	),
						.ra2(	instr[20:16]	),
						.wa3(	writereg	),
						.wd3(	result	),
						.rd1(	srca		),
						.rd2(	writedata      ));

//destination register selection mux						
mux2_5	wrmux(	.in0(	instr[20:16]	),
						.in1(	instr[15:11]	),
						.sel(	regdst			),
						.out(	writereg			));

//register data input selection mux						
mux2_32	resmux(	.in0(	aluresult ),
						.in1(	readdata	),
						.sel(	memtoreg	),
						.out(	result	));
// sign extender to make 32-bit constant						
signext	se(		.a(	instr[15:0]	),
						.y(	signimm		));

/************************************/
/************ ALU Logic **********/
//ALU input B selection mux

mux2_32 srcbmux(	.in0(	writedata ),
						.in1(	signimm 	),
						.sel(	alusrc	),
						.out(	srcb	));
						
//The arithmetic Logic unit
ALU	alu(		.ALUControl( alucontrol	),
					.A( srca 			),
					.B( srcb				),
					.Result(	aluresult		),
					.Zero_Flag(	zero	));
					
/*************************************/

endmodule
